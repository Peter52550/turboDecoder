../../../../lef/BONDPAD.lef