../../../../lef/fsa0m_a_generic_core.lef