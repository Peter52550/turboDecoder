../../../../lef/fsa0m_a_t33_generic_io.lef