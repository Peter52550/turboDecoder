../../../../lef/FSA0M_A_GENERIC_CORE_ANT_V55.lef