../../../../lef/FSA0M_A_T33_GENERIC_IO_ANT_V55.lef