../../../../lef/header6_V55_20ka_cic.lef