module AN2(O, I1, I2);
   output O;
   input I1, I2;
endmodule
module AN2B1(O, I1, B1);
   output O;
   input I1, B1;
endmodule
module AN2B1P(O, I1, B1);
   output O;
   input I1, B1;
endmodule
module AN2B1S(O, I1, B1);
   output O;
   input I1, B1;
endmodule
module AN2B1T(O, I1, B1);
   output O;
   input I1, B1;
endmodule
module AN2P(O, I1, I2);
   output O;
   input I1, I2;
endmodule
module AN2S(O, I1, I2);
   output O;
   input I1, I2;
endmodule
module AN2T(O, I1, I2);
   output O;
   input I1, I2;
endmodule
module AN3(O, I1, I2, I3);
   output O;
   input I1, I2, I3;
endmodule
module AN3B1(O, I1, I2, B1);
   output O;
   input I1, I2, B1;
endmodule
module AN3B1P(O, I1, I2, B1);
   output O;
   input I1, I2, B1;
endmodule
module AN3B1S(O, I1, I2, B1);
   output O;
   input I1, I2, B1;
endmodule
module AN3B1T(O, I1, I2, B1);
   output O;
   input I1, I2, B1;
endmodule
module AN3B2(O, I1, B1, B2);
   output O;
   input I1, B1, B2;
endmodule
module AN3B2P(O, I1, B1, B2);
   output O;
   input I1, B1, B2;
endmodule
module AN3B2S(O, I1, B1, B2);
   output O;
   input I1, B1, B2;
endmodule
module AN3B2T(O, I1, B1, B2);
   output O;
   input I1, B1, B2;
endmodule
module AN3P(O, I1, I2, I3);
   output O;
   input I1, I2, I3;
endmodule
module AN3S(O, I1, I2, I3);
   output O;
   input I1, I2, I3;
endmodule
module AN3T(O, I1, I2, I3);
   output O;
   input I1, I2, I3;
endmodule
module AN4(O, I1, I2, I3, I4);
   output O;
   input I1, I2, I3, I4;
endmodule
module AN4B1(O, I1, I2, I3, B1);
   output O;
   input I1, I2, I3, B1;
endmodule
module AN4B1P(O, I1, I2, I3, B1);
   output O;
   input I1, I2, I3, B1;
endmodule
module AN4B1S(O, I1, I2, I3, B1);
   output O;
   input I1, I2, I3, B1;
endmodule
module AN4B1T(O, I1, I2, I3, B1);
   output O;
   input I1, I2, I3, B1;
endmodule
module AN4P(O, I1, I2, I3, I4);
   output O;
   input I1, I2, I3, I4;
endmodule
module AN4S(O, I1, I2, I3, I4);
   output O;
   input I1, I2, I3, I4;
endmodule
module AN4T(O, I1, I2, I3, I4);
   output O;
   input I1, I2, I3, I4;
endmodule
module ANTENNA(A);
  input A;
endmodule
module AO112(O, A1, B1, C1, C2);
   output O;
   input A1, B1, C1, C2;
endmodule
module AO112P(O, A1, B1, C1, C2);
   output O;
   input A1, B1, C1, C2;
endmodule
module AO112S(O, A1, B1, C1, C2);
   output O;
   input A1, B1, C1, C2;
endmodule
module AO112T(O, A1, B1, C1, C2);
   output O;
   input A1, B1, C1, C2;
endmodule
module AO12(O, A1, B1, B2);
   output O;
   input A1, B1, B2;
endmodule
module AO12P(O, A1, B1, B2);
   output O;
   input A1, B1, B2;
endmodule
module AO12S(O, A1, B1, B2);
   output O;
   input A1, B1, B2;
endmodule
module AO12T(O, A1, B1, B2);
   output O;
   input A1, B1, B2;
endmodule
module AO13(O, A1, B1, B2, B3);
   output O;
   input A1, B1, B2, B3;
endmodule
module AO13P(O, A1, B1, B2, B3);
   output O;
   input A1, B1, B2, B3;
endmodule
module AO13S(O, A1, B1, B2, B3);
   output O;
   input A1, B1, B2, B3;
endmodule
module AO13T(O, A1, B1, B2, B3);
   output O;
   input A1, B1, B2, B3;
endmodule
module AO22(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;
endmodule
module AO222(O, A1, A2, B1, B2, C1, C2);
   output O;
   input A1, A2, B1, B2, C1, C2;
endmodule
module AO222P(O, A1, A2, B1, B2, C1, C2);
   output O;
   input A1, A2, B1, B2, C1, C2;
endmodule
module AO222S(O, A1, A2, B1, B2, C1, C2);
   output O;
   input A1, A2, B1, B2, C1, C2;
endmodule
module AO222T(O, A1, A2, B1, B2, C1, C2);
   output O;
   input A1, A2, B1, B2, C1, C2;
endmodule
module AO22P(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;
endmodule
module AO22S(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;
endmodule
module AO22T(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;
endmodule
module AOI112H(O, A1, B1, C1, C2);
   output O;
   input A1, B1, C1, C2;
endmodule
module AOI112HP(O, A1, B1, C1, C2);
   output O;
   input A1, B1, C1, C2;
endmodule
module AOI112HS(O, A1, B1, C1, C2);
   output O;
   input A1, B1, C1, C2;
endmodule
module AOI112HT(O, A1, B1, C1, C2);
   output O;
   input A1, B1, C1, C2;
endmodule
module AOI12H(O, A1, B1, B2);
   output O;
   input A1, B1, B2;
endmodule
module AOI12HP(O, A1, B1, B2);
   output O;
   input A1, B1, B2;
endmodule
module AOI12HS(O, A1, B1, B2);
   output O;
   input A1, B1, B2;
endmodule
module AOI12HT(O, A1, B1, B2);
   output O;
   input A1, B1, B2;
endmodule
module AOI13H(O, A1, B1, B2, B3);
   output O;
   input A1, B1, B2, B3;
endmodule
module AOI13HP(O, A1, B1, B2, B3);
   output O;
   input A1, B1, B2, B3;
endmodule
module AOI13HS(O, A1, B1, B2, B3);
   output O;
   input A1, B1, B2, B3;
endmodule
module AOI13HT(O, A1, B1, B2, B3);
   output O;
   input A1, B1, B2, B3;
endmodule
module AOI222H(O, A1, A2, B1, B2, C1, C2);
   output O;
   input A1, A2, B1, B2, C1, C2;
endmodule
module AOI222HP(O, A1, A2, B1, B2, C1, C2);
   output O;
   input A1, A2, B1, B2, C1, C2;
endmodule
module AOI222HS(O, A1, A2, B1, B2, C1, C2);
   output O;
   input A1, A2, B1, B2, C1, C2;
endmodule
module AOI22H(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;
endmodule
module AOI22HP(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;
endmodule
module AOI22HT(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;
endmodule
module AOI22S(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;
endmodule
module BHD1(H);
  inout H;
endmodule
module BUF1(O, I);
   output O;
   input I;
endmodule
module BUF12CK(O, I);
   output O;
   input I;
endmodule
module BUF1CK(O, I);
   output O;
   input I;
endmodule
module BUF1S(O, I);
   output O;
   input I;
endmodule
module BUF2(O, I);
   output O;
   input I;
endmodule
module BUF2CK(O, I);
   output O;
   input I;
endmodule
module BUF3(O, I);
   output O;
   input I;
endmodule
module BUF3CK(O, I);
   output O;
   input I;
endmodule
module BUF4(O, I);
   output O;
   input I;
endmodule
module BUF4CK(O, I);
   output O;
   input I;
endmodule
module BUF6(O, I);
   output O;
   input I;
endmodule
module BUF6CK(O, I);
   output O;
   input I;
endmodule
module BUF8(O, I);
   output O;
   input I;
endmodule
module BUF8CK(O, I);
   output O;
   input I;
endmodule
module BUFB1(O, I, EB);
   output O;
   input I, EB;
endmodule
module BUFB2(O, I, EB);
   output O;
   input I, EB;
endmodule
module BUFB3(O, I, EB);
   output O;
   input I, EB;
endmodule
module BUFT1(O, I, E);
   output O;
   input I, E;
endmodule
module BUFT2(O, I, E);
   output O;
   input I, E;
endmodule
module BUFT3(O, I, E);
   output O;
   input I, E;
endmodule
module BUFT4(O, I, E);
   output O;
   input I, E;
endmodule
module CMPE4(OEQ, A0, B0, A1, B1, A2, B2, A3, B3);
   input A0, B0, A1, B1, A2, B2, A3, B3;
   output OEQ;
endmodule
module CMPE4S(OEQ, A0, B0, A1, B1, A2, B2, A3, B3);
   input A0, B0, A1, B1, A2, B2, A3, B3;
   output OEQ;
endmodule
module DBFRBN(Q, QB, D, CKB, RB);
   output Q, QB;
   input D, CKB, RB;
endmodule
module DBFRSBN(Q, QB, D, CKB, RB, SB);
   output Q, QB;
   input D, CKB, RB, SB;
endmodule
module DBHRBN(Q, QB, D, CKB, RB);
   output Q, QB;
   input D, CKB, RB;
endmodule
module DBHRBS(Q, QB, D, CKB, RB);
   output Q, QB;
   input D, CKB, RB;
endmodule
module DBZRBN(Q, QB, D, TD, CKB, SEL, RB);
   output Q, QB;
   input D, CKB, TD, SEL, RB;
endmodule
module DBZRSBN(Q, QB, D, TD, CKB, SEL, RB, SB);
   output Q, QB;
   input D, TD, CKB, RB, SB, SEL;
endmodule
module DELA(O, I);
  output O;
  input I;
endmodule
module DELB(O, I);
  output O;
  input I;
endmodule
module DELC(O, I);
  output O;
  input I;
endmodule
module DFCLRBN(Q, QB, D, CK, RB, LD);
   output Q, QB;
   input D, CK, RB, LD;
endmodule
module DFCRBN(Q, QB, D, CK, RB);
   output Q, QB;
   input D, CK, RB;
endmodule
module DFFN(Q, QB, D, CK);
   output Q, QB;
   input D, CK;
endmodule
module DFFP(Q, QB, D, CK);
   output Q, QB;
   input D, CK;
endmodule
module DFFRBN(Q, QB, D, CK, RB);
   output Q, QB;
   input D, CK, RB;
endmodule
module DFFRBP(Q, QB, D, CK, RB);
   output Q, QB;
   input D, CK, RB;
endmodule
module DFFRBS(Q, QB, D, CK, RB);
   output Q, QB;
   input D, CK, RB;
endmodule
module DFFRBT(Q, QB, D, CK, RB);
   output Q, QB;
   input D, CK, RB;
endmodule
module DFFRSBN(Q, QB, D, CK, RB, SB);
   output Q, QB;
   input D, CK, RB, SB;
endmodule
module DFFS(Q, QB, D, CK);
   output Q, QB;
   input D, CK;
endmodule
module DFFSBN(Q, QB, D, CK, SB);
   output Q, QB;
   input D, CK, SB;
endmodule
module DFTRBN(Q, QZ, D, CK, RB, E);
   output QZ;
   output Q;
   input D,CK, E, RB;
endmodule
module DFTRBS(Q, QZ, D, CK, RB, E);
   output QZ;
   output Q;
   input D,CK, E, RB;
endmodule
module DFZCLRBN(Q, QB, D, TD, CK, RB, SEL, LD);
   output Q, QB;
   input D, TD, CK, RB, SEL, LD;
endmodule
module DFZCRBN(Q, QB, D, TD, CK, SEL, RB);
   output Q, QB;
   input D, TD, CK, SEL, RB;
endmodule
module DFZN(Q, QB, D, TD, CK, SEL);
   output Q, QB;
   input D, CK, TD, SEL;
endmodule
module DFZP(Q, QB, D, TD, CK, SEL);
   output Q, QB;
   input D, CK, TD, SEL;
endmodule
module DFZRBN(Q, QB, D, TD, CK, SEL, RB);
   output Q, QB;
   input D, CK, TD, RB, SEL;
endmodule
module DFZRBP(Q, QB, D, TD, CK, SEL, RB);
   output Q, QB;
   input D, CK, TD, RB, SEL;
endmodule
module DFZRBS(Q, QB, D, TD, CK, SEL, RB);
   output Q, QB;
   input D, CK, TD, RB, SEL;
endmodule
module DFZRBT(Q, QB, D, TD, CK, SEL, RB);
   output Q, QB;
   input D, CK, TD, RB, SEL;
endmodule
module DFZRSBN(Q, QB, D, TD, CK, SEL, RB, SB);
   output Q, QB;
   input D, CK, TD, SB, SEL, RB;
endmodule
module DFZS(Q, QB, D, TD, CK, SEL);
   output Q, QB;
   input D, CK, TD, SEL;
endmodule
module DFZSBN(Q, QB, D, TD, CK, SEL, SB);
   output Q, QB;
   input D, CK, TD, SB, SEL;
endmodule
module DFZTRBN(Q, QZ, D, TD, CK, SEL, RB, E);
   output QZ;
   output Q;
   input D, TD, CK, E, SEL, RB;
endmodule
module DFZTRBS(Q, QZ, D, TD, CK, SEL, RB, E);
   output QZ;
   output Q;
   input D, TD, CK, E, SEL, RB;
endmodule
module DLHN(Q, QB, D, CK);
   output Q, QB;
   input D, CK;
endmodule
module DLHP(Q, QB, D, CK);
   output Q, QB;
   input D, CK;
endmodule
module DLHRBN(Q, QB, D, CK, RB);
   output Q, QB;
   input D, CK, RB;
endmodule
module DLHRBP(Q, QB, D, CK, RB);
   output Q, QB;
   input D, CK, RB;
endmodule
module DLHRBS(Q, QB, D, CK, RB);
   output Q, QB;
   input D, CK, RB;
endmodule
module DLHS(Q, QB, D, CK);
   output Q, QB;
   input D, CK;
endmodule
module FA1(S, CO, A, B, CI);
   output S, CO;
   input A, B, CI;
endmodule
module FA1P(S, CO, A, B, CI);
   output S, CO;
   input A, B, CI;
endmodule
module FA1S(S, CO, A, B, CI);
   output S, CO;
   input A, B, CI;
endmodule
module FA1T(S, CO, A, B, CI);
   output S, CO;
   input A, B, CI;
endmodule
module FA2(S, CO, A, B, CI);
   output S, CO;
   input A, B, CI;
endmodule
module FA2P(S, CO, A, B, CI);
   output S, CO;
   input A, B, CI;
endmodule
module FA2S(S, CO, A, B, CI);
   output S, CO;
   input A, B, CI;
endmodule
module FA3(S, CO, A, B, CI);
   output S, CO;
   input A, B, CI;
endmodule
module FA3P(S, CO, A, B, CI);
   output S, CO;
   input A, B, CI;
endmodule
module FA3S(S, CO, A, B, CI);
   output S, CO;
   input A, B, CI;
endmodule
module FACS1(S, CO0, CO1, A, B, CI0, CI1, CS);
   output S, CO0, CO1;
   input A, B, CI0, CI1, CS;
endmodule
module FACS1P(S, CO0, CO1, A, B, CI0, CI1, CS);
   output S, CO0, CO1;
   input A, B, CI0, CI1, CS;
endmodule
module FACS1S(S, CO0, CO1, A, B, CI0, CI1, CS);
   output S, CO0, CO1;
   input A, B, CI0, CI1, CS;
endmodule
module FACS2(S, CO0, CO1, A, B, CI0, CI1, CS);
   output S, CO0, CO1;
   input A, B, CI0, CI1, CS;
endmodule
module FACS2P(S, CO0, CO1, A, B, CI0, CI1, CS);
   output S, CO0, CO1;
   input A, B, CI0, CI1, CS;
endmodule
module FACS2S(S, CO0, CO1, A, B, CI0, CI1, CS);
   output S, CO0, CO1;
   input A, B, CI0, CI1, CS;
endmodule
module GCKETF(Q, E, TE, CK);
   output Q;
   input E, TE, CK;
endmodule
module GCKETN(Q, E, TE, CK);
   output Q;
   input E, TE, CK;
endmodule
module GCKETP(Q, E, TE, CK);
   output Q;
   input E, TE, CK;
endmodule
module GCKETT(Q, E, TE, CK);
   output Q;
   input E, TE, CK;
endmodule
module HA1(S, C, A, B);
   output S, C;
   input A, B;
endmodule
module HA1P(S, C, A, B);
   output S, C;
   input A, B;
endmodule
module HA1S(S, C, A, B);
   output S, C;
   input A, B;
endmodule
module HA1T(S, C, A, B);
   output S, C;
   input A, B;
endmodule
module HA2(S, C, A, B);
   output S, C;
   input A, B;
endmodule
module HA2P(S, C, A, B);
   output S, C;
   input A, B;
endmodule
module HA2T(S, C, A, B);
   output S, C;
   input A, B;
endmodule
module HA3(S, C, A, B);
   output S, C;
   input A, B;
endmodule
module HA3P(S, C, A, B);
   output S, C;
   input A, B;
endmodule
module HA3T(S, C, A, B);
   output S, C;
   input A, B;
endmodule
module INV1(O, I);
   output O;
   input I;
endmodule
module INV12(O, I);
   output O;
   input I;
endmodule
module INV12CK(O, I);
   output O;
   input I;
endmodule
module INV1CK(O, I);
   output O;
   input I;
endmodule
module INV1S(O, I);
   output O;
   input I;
endmodule
module INV2(O, I);
   output O;
   input I;
endmodule
module INV2CK(O, I);
   output O;
   input I;
endmodule
module INV3(O, I);
   output O;
   input I;
endmodule
module INV3CK(O, I);
   output O;
   input I;
endmodule
module INV4(O, I);
   output O;
   input I;
endmodule
module INV4CK(O, I);
   output O;
   input I;
endmodule
module INV6(O, I);
   output O;
   input I;
endmodule
module INV6CK(O, I);
   output O;
   input I;
endmodule
module INV8(O, I);
   output O;
   input I;
endmodule
module INV8CK(O, I);
   output O;
   input I;
endmodule
module INVT1(O, I, E);
   output O;
   input I, E;
endmodule
module INVT2(O, I, E);
   output O;
   input I, E;
endmodule
module INVT4(O, I, E);
   output O;
   input I, E;
endmodule
module JKFN(Q, QB, J, K, CK);
   output Q, QB;
   input J, K, CK;
endmodule
module JKFRBN(Q, QB, J, K, CK, RB);
   output Q, QB;
   input J, K, CK, RB;
endmodule
module JKFRBP(Q, QB, J, K, CK, RB);
   output Q, QB;
   input J, K, CK, RB;
endmodule
module JKZN(Q, QB, J, K, TD, CK, SEL);
   output Q, QB;
   input J, K, CK, TD, SEL;
endmodule
module JKZRBN(Q, QB, J, K, TD, CK, SEL, RB);
   output Q, QB;
   input J, K, CK, TD, SEL, RB;
endmodule
module JKZRBP(Q, QB, J, K, TD, CK, SEL, RB);
   output Q, QB;
   input J, K, CK, TD, SEL, RB;
endmodule
module MAO222(O, A1, B1, C1);
   output O;
   input A1, B1, C1;
endmodule
module MAO222P(O, A1, B1, C1);
   output O;
   input A1, B1, C1;
endmodule
module MAO222S(O, A1, B1, C1);
   output O;
   input A1, B1, C1;
endmodule
module MAO222T(O, A1, B1, C1);
   output O;
   input A1, B1, C1;
endmodule
module MAOI1(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;
endmodule
module MAOI1H(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;
endmodule
module MAOI1HP(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;
endmodule
module MAOI1HT(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;
endmodule
module MAOI1S(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;
endmodule
module MOAI1(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;
endmodule
module MOAI1H(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;
endmodule
module MOAI1HP(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;
endmodule
module MOAI1HT(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;
endmodule
module MOAI1S(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;
endmodule
module MULBE(S, M, Z, M0, M1, M2);
   output S, M, Z;
   input M0, M1, M2;
endmodule
module MULBEP(S, M, Z, M0, M1, M2);
   output S, M, Z;
   input M0, M1, M2;
endmodule
module MULBET(S, M, Z, M0, M1, M2);
   output S, M, Z;
   input M0, M1, M2;
endmodule
module MULPA(P, S, M, Z, M0, M1);
   output P;
   input S, M, Z, M1, M0;
endmodule
module MULPAP(P, S, M, Z, M0, M1);
   output P;
   input S, M, Z, M1, M0;
endmodule
module MULPAT(P, S, M, Z, M0, M1);
   output P;
   input S, M, Z, M1, M0;
endmodule
module MUX2(O, S, A, B);
   input A, B, S;
   output O;
endmodule
module MUX2F(O, S, A, B);
   input A, B, S;
   output O;
endmodule
module MUX2P(O, S, A, B);
   input A, B, S;
   output O;
endmodule
module MUX2S(O, S, A, B);
   input A, B, S;
   output O;
endmodule
module MUX2T(O, S, A, B);
   input A, B, S;
   output O;
endmodule
module MUX3(O, S0, S1, A, B, C);
   input A, B, C, S0, S1;
   output O;
endmodule
module MUX3P(O, S0, S1, A, B, C);
   input A, B, C, S0, S1;
   output O;
endmodule
module MUX3S(O, S0, S1, A, B, C);
   input A, B, C, S0, S1;
   output O;
endmodule
module MUX3T(O, S0, S1, A, B, C);
   input A, B, C, S0, S1;
   output O;
endmodule
module MUX4(O, S0, S1, A, B, C, D);
   output O;
   input S0, S1, A, B, C, D;
endmodule
module MUX4P(O, S0, S1, A, B, C, D);
   output O;
   input S0, S1, A, B, C, D;
endmodule
module MUX4S(O, S0, S1, A, B, C, D);
   output O;
   input S0, S1, A, B, C, D;
endmodule
module MUX4T(O, S0, S1, A, B, C, D);
   output O;
   input S0, S1, A, B, C, D;
endmodule
module MUXB2(O, S, A, B, EB);
   input A, B, S, EB;
   output O;
endmodule
module MUXB2P(O, S, A, B, EB);
   input A, B, S, EB;
   output O;
endmodule
module MUXB2S(O, S, A, B, EB);
   input A, B, S, EB;
   output O;
endmodule
module MUXB2T(O, S, A, B, EB);
   input A, B, S, EB;
   output O;
endmodule
module MUXB4(O, S0, S1, A, B, C, D, EB);
   output O;
   input S0, S1, A, B, C, D, EB;
endmodule
module MUXB4P(O, S0, S1, A, B, C, D, EB);
   output O;
   input S0, S1, A, B, C, D, EB;
endmodule
module MUXB4S(O, S0, S1, A, B, C, D, EB);
   output O;
   input S0, S1, A, B, C, D, EB;
endmodule
module MUXB4T(O, S0, S1, A, B, C, D, EB);
   output O;
   input S0, S1, A, B, C, D, EB;
endmodule
module MXL2H(OB, S, A, B);
   input A, B, S;
   output OB;
endmodule
module MXL2HF(OB, S, A, B);
   input A, B, S;
   output OB;
endmodule
module MXL2HP(OB, S, A, B);
   input A, B, S;
   output OB;
endmodule
module MXL2HS(OB, S, A, B);
   input A, B, S;
   output OB;
endmodule
module MXL2HT(OB, S, A, B);
   input A, B, S;
   output OB;
endmodule
module MXL3(OB, S0, S1, A, B, C);
   input A, B, C, S0, S1;
   output OB;
endmodule
module MXL3P(OB, S0, S1, A, B, C);
   input A, B, C, S0, S1;
   output OB;
endmodule
module MXL3S(OB, S0, S1, A, B, C);
   input A, B, C, S0, S1;
   output OB;
endmodule
module MXL3T(OB, S0, S1, A, B, C);
   input A, B, C, S0, S1;
   output OB;
endmodule
module ND2(O, I1, I2);
   output O;
   input I1, I2;
endmodule
module ND2F(O, I1, I2);
   output O;
   input I1, I2;
endmodule
module ND2P(O, I1, I2);
   output O;
   input I1, I2;
endmodule
module ND2S(O, I1, I2);
   output O;
   input I1, I2;
endmodule
module ND2T(O, I1, I2);
   output O;
   input I1, I2;
endmodule
module ND3(O, I1, I2, I3);
   output O;
   input I1, I2, I3;
endmodule
module ND3HT(O, I1, I2, I3);
   output O;
   input I1, I2, I3;
endmodule
module ND3P(O, I1, I2, I3);
   output O;
   input I1, I2, I3;
endmodule
module ND3S(O, I1, I2, I3);
   output O;
   input I1, I2, I3;
endmodule
module ND4(O, I1, I2, I3, I4);
   output O;
   input I1, I2, I3, I4;
endmodule
module ND4P(O, I1, I2, I3, I4);
   output O;
   input I1, I2, I3, I4;
endmodule
module ND4S(O, I1, I2, I3, I4);
   output O;
   input I1, I2, I3, I4;
endmodule
module ND4T(O, I1, I2, I3, I4);
   output O;
   input I1, I2, I3, I4;
endmodule
module NR2(O, I1, I2);
   output O;
   input I1, I2;
endmodule
module NR2F(O, I1, I2);
   output O;
   input I1, I2;
endmodule
module NR2P(O, I1, I2);
   output O;
   input I1, I2;
endmodule
module NR2T(O, I1, I2);
   output O;
   input I1, I2;
endmodule
module NR3(O, I1, I2, I3);
   output O;
   input I1, I2, I3;
endmodule
module NR3H(O, I1, I2, I3);
   output O;
   input I1, I2, I3;
endmodule
module NR3HP(O, I1, I2, I3);
   output O;
   input I1, I2, I3;
endmodule
module NR3HT(O, I1, I2, I3);
   output O;
   input I1, I2, I3;
endmodule
module NR4(O, I1, I2, I3, I4);
   output O;
   input I1, I2, I3, I4;
endmodule
module NR4P(O, I1, I2, I3, I4);
   output O;
   input I1, I2, I3, I4;
endmodule
module NR4S(O, I1, I2, I3, I4);
   output O;
   input I1, I2, I3, I4;
endmodule
module NR4T(O, I1, I2, I3, I4);
   output O;
   input I1, I2, I3, I4;
endmodule
module OA112(O, A1, B1, C1, C2);
   output O;
   input A1, B1, C1, C2;
endmodule
module OA112P(O, A1, B1, C1, C2);
   output O;
   input A1, B1, C1, C2;
endmodule
module OA112S(O, A1, B1, C1, C2);
   output O;
   input A1, B1, C1, C2;
endmodule
module OA112T(O, A1, B1, C1, C2);
   output O;
   input A1, B1, C1, C2;
endmodule
module OA12(O, A1, B1, B2);
   output O;
   input A1, B1, B2;
endmodule
module OA12P(O, A1, B1, B2);
   output O;
   input A1, B1, B2;
endmodule
module OA12S(O, A1, B1, B2);
   output O;
   input A1, B1, B2;
endmodule
module OA12T(O, A1, B1, B2);
   output O;
   input A1, B1, B2;
endmodule
module OA13(O, A1, B1, B2, B3);
   output O;
   input A1, B1, B2, B3;
endmodule
module OA13P(O, A1, B1, B2, B3);
   output O;
   input A1, B1, B2, B3;
endmodule
module OA13S(O, A1, B1, B2, B3);
   output O;
   input A1, B1, B2, B3;
endmodule
module OA13T(O, A1, B1, B2, B3);
   output O;
   input A1, B1, B2, B3;
endmodule
module OA22(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;
endmodule
module OA222(O, A1, A2, B1, B2, C1, C2);
   output O;
   input A1, A2, B1, B2, C1, C2;
endmodule
module OA222P(O, A1, A2, B1, B2, C1, C2);
   output O;
   input A1, A2, B1, B2, C1, C2;
endmodule
module OA222S(O, A1, A2, B1, B2, C1, C2);
   output O;
   input A1, A2, B1, B2, C1, C2;
endmodule
module OA222T(O, A1, A2, B1, B2, C1, C2);
   output O;
   input A1, A2, B1, B2, C1, C2;
endmodule
module OA22P(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;
endmodule
module OA22S(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;
endmodule
module OA22T(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;
endmodule
module OAI112H(O, A1, B1, C1, C2);
   output O;
   input A1, B1, C1, C2;
endmodule
module OAI112HP(O, A1, B1, C1, C2);
   output O;
   input A1, B1, C1, C2;
endmodule
module OAI112HS(O, A1, B1, C1, C2);
   output O;
   input A1, B1, C1, C2;
endmodule
module OAI112HT(O, A1, B1, C1, C2);
   output O;
   input A1, B1, C1, C2;
endmodule
module OAI12H(O, A1, B1, B2);
   output O;
   input A1, B1, B2;
endmodule
module OAI12HP(O, A1, B1, B2);
   output O;
   input A1, B1, B2;
endmodule
module OAI12HS(O, A1, B1, B2);
   output O;
   input A1, B1, B2;
endmodule
module OAI12HT(O, A1, B1, B2);
   output O;
   input A1, B1, B2;
endmodule
module OAI13H(O, A1, B1, B2, B3);
   output O;
   input A1, B1, B2, B3;
endmodule
module OAI13HP(O, A1, B1, B2, B3);
   output O;
   input A1, B1, B2, B3;
endmodule
module OAI13HS(O, A1, B1, B2, B3);
   output O;
   input A1, B1, B2, B3;
endmodule
module OAI13HT(O, A1, B1, B2, B3);
   output O;
   input A1, B1, B2, B3;
endmodule
module OAI222H(O, A1, A2, B1, B2, C1, C2);
   output O;
   input A1, A2, B1, B2, C1, C2;
endmodule
module OAI222HP(O, A1, A2, B1, B2, C1, C2);
   output O;
   input A1, A2, B1, B2, C1, C2;
endmodule
module OAI222HT(O, A1, A2, B1, B2, C1, C2);
   output O;
   input A1, A2, B1, B2, C1, C2;
endmodule
module OAI222S(O, A1, A2, B1, B2, C1, C2);
   output O;
   input A1, A2, B1, B2, C1, C2;
endmodule
module OAI22H(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;
endmodule
module OAI22HP(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;
endmodule
module OAI22HT(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;
endmodule
module OAI22S(O, A1, A2, B1, B2);
   output O;
   input A1, A2, B1, B2;
endmodule
module OR2(O, I1, I2);
   output O;
   input I1, I2;
endmodule
module OR2B1(O, I1, B1);
   output O;
   input I1, B1;
endmodule
module OR2B1P(O, I1, B1);
   output O;
   input I1, B1;
endmodule
module OR2B1S(O, I1, B1);
   output O;
   input I1, B1;
endmodule
module OR2B1T(O, I1, B1);
   output O;
   input I1, B1;
endmodule
module OR2P(O, I1, I2);
   output O;
   input I1, I2;
endmodule
module OR2S(O, I1, I2);
   output O;
   input I1, I2;
endmodule
module OR2T(O, I1, I2);
   output O;
   input I1, I2;
endmodule
module OR3(O, I1, I2, I3);
   output O;
   input I1, I2, I3;
endmodule
module OR3B1(O, I1, I2, B1);
   output O;
   input I1, I2, B1;
endmodule
module OR3B1P(O, I1, I2, B1);
   output O;
   input I1, I2, B1;
endmodule
module OR3B1S(O, I1, I2, B1);
   output O;
   input I1, I2, B1;
endmodule
module OR3B1T(O, I1, I2, B1);
   output O;
   input I1, I2, B1;
endmodule
module OR3B2(O, I1, B1, B2);
   output O;
   input I1, B1, B2;
endmodule
module OR3B2P(O, I1, B1, B2);
   output O;
   input I1, B1, B2;
endmodule
module OR3B2S(O, I1, B1, B2);
   output O;
   input I1, B1, B2;
endmodule
module OR3B2T(O, I1, B1, B2);
   output O;
   input I1, B1, B2;
endmodule
module OR3P(O, I1, I2, I3);
   output O;
   input I1, I2, I3;
endmodule
module OR3S(O, I1, I2, I3);
   output O;
   input I1, I2, I3;
endmodule
module OR3T(O, I1, I2, I3);
   output O;
   input I1, I2, I3;
endmodule
module PDI(O, EB);
   input EB;
   output O;
endmodule
module PDIX(O, EB);
   input EB;
   output O;
endmodule
module PUI(O, E);
   input E;
   output O;
endmodule
module QDBHN(Q, D, CKB);
   output Q;
   input D, CKB;
endmodule
module QDBHS(Q, D, CKB);
   output Q;
   input D, CKB;
endmodule
module QDFFN(Q, D, CK);
   output Q;
   input D, CK;
endmodule
module QDFFP(Q, D, CK);
   output Q;
   input D, CK;
endmodule
module QDFFRBN(Q, D, CK, RB);
   output Q;
   input D, CK, RB;
endmodule
module QDFFRBP(Q, D, CK, RB);
   output Q;
   input D, CK, RB;
endmodule
module QDFFRBS(Q, D, CK, RB);
   output Q;
   input D, CK, RB;
endmodule
module QDFFRBT(Q, D, CK, RB);
   output Q;
   input D, CK, RB;
endmodule
module QDFFRSBN(Q, D, CK, RB, SB);
   output Q;
   input D, CK, RB, SB;
endmodule
module QDFFS(Q, D, CK);
   output Q;
   input D, CK;
endmodule
module QDFZN(Q, D, TD, CK, SEL);
   output Q;
   input D, CK, TD, SEL;
endmodule
module QDFZP(Q, D, TD, CK, SEL);
   output Q;
   input D, CK, TD, SEL;
endmodule
module QDFZRBN(Q, D, TD, CK, SEL, RB);
   output Q;
   input D, CK, TD, RB, SEL;
endmodule
module QDFZRBP(Q, D, TD, CK, SEL, RB);
   output Q;
   input D, CK, TD, RB, SEL;
endmodule
module QDFZRBS(Q, D, TD, CK, SEL, RB);
   output Q;
   input D, CK, TD, RB, SEL;
endmodule
module QDFZRBT(Q, D, TD, CK, SEL, RB);
   output Q;
   input D, CK, TD, RB, SEL;
endmodule
module QDFZRSBN(Q, D, TD, CK, SEL, RB, SB);
   output Q;
   input D, TD, CK, RB, SB, SEL;
endmodule
module QDFZS(Q, D, TD, CK, SEL);
   output Q;
   input D, CK, TD, SEL;
endmodule
module QDLHN(Q, D, CK);
   output Q;
   input D, CK;
endmodule
module QDLHP(Q, D, CK);
   output Q;
   input D, CK;
endmodule
module QDLHRBN(Q, D, CK, RB);
   output Q;
   input D, CK, RB;
endmodule
module QDLHRBP(Q, D, CK, RB);
   output Q;
   input D, CK, RB;
endmodule
module QDLHRBS(Q, D, CK, RB);
   output Q;
   input D, CK, RB;
endmodule
module QDLHS(Q, D, CK);
   output Q;
   input D, CK;
endmodule
module QDLHSN(Q, D, CK, S);
   input D, CK, S;
   output Q;
endmodule
module RAM2(QB, QBZ, D, W, RD);
   output QBZ;
   input D, W, RD;
   output QB;
endmodule
module RAM2S(QB, QBZ, D, W, RD);
   output QBZ;
   input D, W, RD;
   output QB;
endmodule
module RAM3(Q, QZ, D, W, RD);
   output QZ;
   input D, W, RD;
   output Q;
endmodule
module RAM3S(Q, QZ, D, W, RD);
   output QZ;
   input D, W, RD;
   output Q;
endmodule
module RAM5(QZ0, QZ1, D, W, RD0, RD1);
   output QZ0, QZ1;
   input D, W, RD0, RD1;
endmodule
module RAM5S(QZ0, QZ1, D, W, RD0, RD1);
   output QZ0, QZ1;
   input D, W, RD0, RD1;
endmodule
module TIE0(O);
  output O;
endmodule
module TIE1(O);
  output O;
endmodule
module XNR2H(O, I1, I2);
   output O;
   input I1, I2;
endmodule
module XNR2HP(O, I1, I2);
   output O;
   input I1, I2;
endmodule
module XNR2HS(O, I1, I2);
   output O;
   input I1, I2;
endmodule
module XNR2HT(O, I1, I2);
   output O;
   input I1, I2;
endmodule
module XNR3(O, I1, I2, I3);
   output O;
   input I1, I2, I3;
endmodule
module XNR3P(O, I1, I2, I3);
   output O;
   input I1, I2, I3;
endmodule
module XNR3S(O, I1, I2, I3);
   output O;
   input I1, I2, I3;
endmodule
module XNR3T(O, I1, I2, I3);
   output O;
   input I1, I2, I3;
endmodule
module XNR4(O, I1, I2, I3, I4);
   output O;
   input I1, I2, I3, I4;
endmodule
module XNR4P(O, I1, I2, I3, I4);
   output O;
   input I1, I2, I3, I4;
endmodule
module XNR4S(O, I1, I2, I3, I4);
   output O;
   input I1, I2, I3, I4;
endmodule
module XNR4T(O, I1, I2, I3, I4);
   output O;
   input I1, I2, I3, I4;
endmodule
module XOR2H(O, I1, I2);
   output O;
   input I1, I2;
endmodule
module XOR2HP(O, I1, I2);
   output O;
   input I1, I2;
endmodule
module XOR2HS(O, I1, I2);
   output O;
   input I1, I2;
endmodule
module XOR2HT(O, I1, I2);
   output O;
   input I1, I2;
endmodule
module XOR3(O, I1, I2, I3);
   output O;
   input I1, I2, I3;
endmodule
module XOR3P(O, I1, I2, I3);
   output O;
   input I1, I2, I3;
endmodule
module XOR3S(O, I1, I2, I3);
   output O;
   input I1, I2, I3;
endmodule
module XOR3T(O, I1, I2, I3);
   output O;
   input I1, I2, I3;
endmodule
module XOR4(O, I1, I2, I3, I4);
   output O;
   input I1, I2, I3, I4;
endmodule
module XOR4P(O, I1, I2, I3, I4);
   output O;
   input I1, I2, I3, I4;
endmodule
module XOR4S(O, I1, I2, I3, I4);
   output O;
   input I1, I2, I3, I4;
endmodule
module XOR4T(O, I1, I2, I3, I4);
   output O;
   input I1, I2, I3, I4;
endmodule
