* SPICE NETLIST
***************************************

.SUBCKT L POS NEG SUB
.ENDS
***************************************
.SUBCKT ICV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT YA2GSC O E E2 E8 E4 I SR
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_2 1 2 3 4 5 6 7
** N=7 EP=7 IP=16 FDC=0
X0 5 1 2 2 2 3 2 YA2GSC $T=1080850 752120 0 90 $X=845870 $Y=754030
X1 6 1 2 2 2 4 2 YA2GSC $T=1080850 813300 0 90 $X=845870 $Y=815210
.ENDS
***************************************
.SUBCKT ICV_3 1 2 3 4 5
** N=5 EP=5 IP=8 FDC=0
X0 4 1 2 2 2 3 2 YA2GSC $T=1080850 690940 0 90 $X=845870 $Y=692850
.ENDS
***************************************
.SUBCKT ICV_4 2 3 4 5 10
** N=10 EP=5 IP=8 FDC=0
X0 2 3 4 4 4 5 4 YA2GSC $T=1080850 629760 0 90 $X=845870 $Y=631670
.ENDS
***************************************
.SUBCKT ICV_5 1 2 3 5 10
** N=15 EP=5 IP=8 FDC=0
X0 5 1 2 2 2 3 2 YA2GSC $T=1080850 446220 0 90 $X=845870 $Y=448130
.ENDS
***************************************
.SUBCKT ICV_6 1 2 3 4 5
** N=5 EP=5 IP=8 FDC=0
X0 4 1 2 2 2 3 2 YA2GSC $T=1080850 385040 0 90 $X=845870 $Y=386950
.ENDS
***************************************
.SUBCKT ICV_7 1 2 3 4 5 6 7
** N=7 EP=7 IP=16 FDC=0
X0 5 1 2 2 2 3 2 YA2GSC $T=1080850 262680 0 90 $X=845870 $Y=264590
X1 6 1 2 2 2 4 2 YA2GSC $T=1080850 323860 0 90 $X=845870 $Y=325770
.ENDS
***************************************
.SUBCKT ICV_8
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT XMC SMT I PU PD O
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_9 1 2 3 4 5 6
** N=6 EP=6 IP=12 FDC=0
X0 1 3 1 1 2 XMC $T=1110080 -829830 0 90 $X=875100 $Y=-827980
X1 1 5 1 1 4 XMC $T=1110080 -780310 0 90 $X=875100 $Y=-778460
.ENDS
***************************************
.SUBCKT ICV_10
** N=9 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_11
** N=8 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_12
** N=6 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_13
** N=8 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT BUF2CK I O GND VCC
** N=6 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_14 1 2 3 4 9
** N=9 EP=5 IP=5 FDC=0
X0 1 2 4 3 BUF2CK $T=730360 441840 1 0 $X=730360 $Y=436420
.ENDS
***************************************
.SUBCKT ICV_15
** N=10 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_16 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=16 FDC=0
X0 1 2 3 3 4 5 4 YA2GSC $T=0 -786720 0 270 $X=0 $Y=-819590
X1 6 2 3 3 3 7 3 YA2GSC $T=0 -728200 0 270 $X=0 $Y=-761070
.ENDS
***************************************
.SUBCKT ICV_17 5 6 7 8 9 10 11 30
** N=40 EP=8 IP=18 FDC=0
X0 5 7 5 5 6 XMC $T=631750 1110080 0 180 $X=599560 $Y=875100
X1 5 9 5 5 8 XMC $T=681270 1110080 0 180 $X=649080 $Y=875100
X2 5 11 5 5 10 XMC $T=730790 1110080 0 180 $X=698600 $Y=875100
.ENDS
***************************************
.SUBCKT ICV_18
** N=29 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT TIE0 O VCC GND
** N=5 EP=3 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT QDFFRBT D CK RB GND VCC Q
** N=17 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT QDFFRBN D CK RB VCC GND Q
** N=18 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_19 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 17 18 19 20 22
** N=22 EP=20 IP=53 FDC=0
X0 8 19 20 TIE0 $T=562340 673680 0 0 $X=562340 $Y=673300
X1 12 4 3 20 19 15 QDFFRBT $T=591480 693840 1 0 $X=591480 $Y=688420
X2 18 4 3 20 19 13 QDFFRBT $T=610080 703920 1 180 $X=596440 $Y=703540
X3 6 4 3 19 20 1 QDFFRBN $T=551800 693840 1 180 $X=540020 $Y=693460
X4 5 4 3 19 20 2 QDFFRBN $T=552420 703920 1 180 $X=540640 $Y=703540
X5 9 4 3 19 20 7 QDFFRBN $T=564820 703920 1 180 $X=553040 $Y=703540
X6 11 4 3 19 20 10 QDFFRBN $T=582800 703920 0 180 $X=571020 $Y=698500
X7 17 4 3 19 20 14 QDFFRBN $T=613180 693840 1 180 $X=601400 $Y=693460
.ENDS
***************************************
.SUBCKT FA1S CO VCC A B CI GND S
** N=14 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NR2 I1 VCC O I2 GND
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT HA1 A B C GND VCC S
** N=12 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INV1S I VCC O GND
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_20 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 58
** N=163 EP=54 IP=619 FDC=0
X0 52 47 48 19 11 46 QDFFRBT $T=607600 633360 1 180 $X=593960 $Y=632980
X1 45 47 48 19 11 50 QDFFRBT $T=594580 653520 0 0 $X=594580 $Y=653140
X2 70 11 75 85 69 19 8 FA1S $T=502200 643440 1 180 $X=490420 $Y=643060
X3 67 11 63 73 60 19 14 FA1S $T=491660 593040 0 0 $X=491660 $Y=592660
X4 68 11 64 62 77 19 74 FA1S $T=491660 623280 0 0 $X=491660 $Y=622900
X5 72 11 76 78 74 19 65 FA1S $T=504060 613200 1 180 $X=492280 $Y=612820
X6 71 11 67 65 15 19 25 FA1S $T=493520 603120 1 0 $X=493520 $Y=597700
X7 75 11 68 88 79 19 66 FA1S $T=507780 633360 1 180 $X=496000 $Y=632980
X8 69 11 72 66 71 19 18 FA1S $T=499100 633360 1 0 $X=499100 $Y=627940
X9 90 11 86 81 89 19 79 FA1S $T=514600 643440 0 0 $X=514600 $Y=643060
X10 95 11 92 93 87 19 88 FA1S $T=520180 633360 0 0 $X=520180 $Y=632980
X11 101 11 100 99 103 19 110 FA1S $T=527000 623280 0 0 $X=527000 $Y=622900
X12 102 11 97 98 91 19 107 FA1S $T=527620 633360 1 0 $X=527620 $Y=627940
X13 104 11 90 107 105 19 85 FA1S $T=539400 643440 1 180 $X=527620 $Y=643060
X14 120 11 121 95 110 19 105 FA1S $T=552420 633360 1 180 $X=540640 $Y=632980
X15 116 11 104 122 70 19 34 FA1S $T=540640 643440 0 0 $X=540640 $Y=643060
X16 32 11 113 111 114 19 124 FA1S $T=541880 593040 0 0 $X=541880 $Y=592660
X17 119 11 109 115 106 19 125 FA1S $T=543120 613200 1 0 $X=543120 $Y=607780
X18 128 11 118 132 101 19 140 FA1S $T=550560 623280 0 0 $X=550560 $Y=622900
X19 129 11 136 125 102 19 138 FA1S $T=551800 633360 1 0 $X=551800 $Y=627940
X20 133 11 120 140 138 19 122 FA1S $T=564820 633360 1 180 $X=553040 $Y=632980
X21 131 11 137 123 108 19 147 FA1S $T=553660 593040 0 0 $X=553660 $Y=592660
X22 145 11 143 141 135 19 152 FA1S $T=565440 613200 0 0 $X=565440 $Y=612820
X23 146 11 144 134 139 19 136 FA1S $T=566680 623280 0 0 $X=566680 $Y=622900
X24 151 11 149 119 146 19 158 FA1S $T=572880 623280 1 0 $X=572880 $Y=617860
X25 38 11 124 145 151 19 160 FA1S $T=575980 603120 0 0 $X=575980 $Y=602740
X26 153 11 147 152 128 19 159 FA1S $T=575980 613200 1 0 $X=575980 $Y=607780
X27 156 11 158 129 159 19 150 FA1S $T=588380 633360 0 180 $X=576600 $Y=627940
X28 40 11 39 36 155 19 44 FA1S $T=577840 593040 1 0 $X=577840 $Y=587620
X29 155 11 148 131 41 19 162 FA1S $T=577840 603120 1 0 $X=577840 $Y=597700
X30 157 11 156 161 154 19 42 FA1S $T=578460 613200 0 0 $X=578460 $Y=612820
X31 154 11 133 150 116 19 43 FA1S $T=578460 633360 0 0 $X=578460 $Y=632980
X32 163 11 162 153 160 19 161 FA1S $T=590860 603120 0 0 $X=590860 $Y=602740
X33 51 11 163 49 157 19 53 FA1S $T=603260 593040 1 0 $X=603260 $Y=587620
X34 1 11 59 2 19 NR2 $T=481120 593040 0 0 $X=481120 $Y=592660
X35 4 11 6 61 19 NR2 $T=485460 603120 0 0 $X=485460 $Y=602740
X36 2 11 62 61 19 NR2 $T=489180 613200 0 0 $X=489180 $Y=612820
X37 1 11 63 10 19 NR2 $T=490420 593040 1 0 $X=490420 $Y=587620
X38 1 11 64 12 19 NR2 $T=492280 613200 1 0 $X=492280 $Y=607780
X39 2 11 73 17 19 NR2 $T=509020 593040 0 0 $X=509020 $Y=592660
X40 10 11 77 17 19 NR2 $T=509020 623280 0 0 $X=509020 $Y=622900
X41 10 11 87 61 19 NR2 $T=514600 633360 1 0 $X=514600 $Y=627940
X42 21 11 80 61 19 NR2 $T=515220 613200 1 0 $X=515220 $Y=607780
X43 12 11 86 17 19 NR2 $T=515220 623280 0 0 $X=515220 $Y=622900
X44 4 11 83 22 19 NR2 $T=516460 603120 0 0 $X=516460 $Y=602740
X45 2 11 93 22 19 NR2 $T=518940 623280 0 0 $X=518940 $Y=622900
X46 1 11 92 23 19 NR2 $T=519560 613200 1 0 $X=519560 $Y=607780
X47 21 11 82 22 19 NR2 $T=519560 613200 0 0 $X=519560 $Y=612820
X48 4 11 84 27 19 NR2 $T=522660 603120 0 0 $X=522660 $Y=602740
X49 12 11 97 61 19 NR2 $T=523280 623280 0 0 $X=523280 $Y=622900
X50 21 11 94 27 19 NR2 $T=523900 613200 1 0 $X=523900 $Y=607780
X51 1 11 109 26 19 NR2 $T=526380 603120 0 180 $X=524520 $Y=597700
X52 10 11 98 22 19 NR2 $T=524520 623280 1 0 $X=524520 $Y=617860
X53 21 11 16 17 19 NR2 $T=525760 593040 1 0 $X=525760 $Y=587620
X54 2 11 99 27 19 NR2 $T=528240 613200 1 0 $X=528240 $Y=607780
X55 1 11 100 29 19 NR2 $T=529480 603120 0 0 $X=529480 $Y=602740
X56 23 11 103 17 19 NR2 $T=532580 613200 1 0 $X=532580 $Y=607780
X57 4 11 96 30 19 NR2 $T=532580 613200 0 0 $X=532580 $Y=612820
X58 26 11 108 17 19 NR2 $T=535680 593040 0 0 $X=535680 $Y=592660
X59 26 11 113 61 19 NR2 $T=535680 603120 0 0 $X=535680 $Y=602740
X60 29 11 106 17 19 NR2 $T=538780 613200 0 180 $X=536920 $Y=607780
X61 31 11 111 2 19 NR2 $T=540020 593040 0 0 $X=540020 $Y=592660
X62 21 11 117 30 19 NR2 $T=542500 613200 0 0 $X=542500 $Y=612820
X63 10 11 114 33 19 NR2 $T=543120 593040 1 0 $X=543120 $Y=587620
X64 2 11 115 30 19 NR2 $T=543120 603120 0 0 $X=543120 $Y=602740
X65 4 11 112 33 19 NR2 $T=543120 623280 0 0 $X=543120 $Y=622900
X66 2 11 130 33 19 NR2 $T=545600 603120 1 0 $X=545600 $Y=597700
X67 21 11 126 33 19 NR2 $T=550560 613200 1 180 $X=548700 $Y=612820
X68 10 11 123 30 19 NR2 $T=553660 593040 0 180 $X=551800 $Y=587620
X69 4 11 127 31 19 NR2 $T=551800 603120 0 0 $X=551800 $Y=602740
X70 31 11 142 21 19 NR2 $T=559860 603120 0 180 $X=558000 $Y=597700
X71 12 11 137 27 19 NR2 $T=559860 593040 1 0 $X=559860 $Y=587620
X72 12 11 139 22 19 NR2 $T=559860 603120 0 0 $X=559860 $Y=602740
X73 10 11 134 27 19 NR2 $T=560480 613200 1 0 $X=560480 $Y=607780
X74 23 11 141 22 19 NR2 $T=566060 593040 1 0 $X=566060 $Y=587620
X75 23 11 144 61 19 NR2 $T=567920 603120 0 0 $X=567920 $Y=602740
X76 29 11 143 61 19 NR2 $T=567920 613200 1 0 $X=567920 $Y=607780
X77 29 11 35 22 19 NR2 $T=571640 593040 0 180 $X=569780 $Y=587620
X78 23 11 37 27 19 NR2 $T=574120 593040 1 0 $X=574120 $Y=587620
X79 59 16 60 19 11 5 HA1 $T=478640 593040 1 0 $X=478640 $Y=587620
X80 80 83 76 19 11 13 HA1 $T=510260 613200 0 180 $X=502200 $Y=607780
X81 82 84 81 19 11 78 HA1 $T=513360 613200 1 180 $X=505300 $Y=612820
X82 94 96 91 19 11 89 HA1 $T=526380 633360 0 180 $X=518320 $Y=627940
X83 117 112 118 19 11 121 HA1 $T=541260 633360 1 0 $X=541260 $Y=627940
X84 126 127 135 19 11 132 HA1 $T=554900 613200 0 0 $X=554900 $Y=612820
X85 130 142 148 19 11 149 HA1 $T=566680 603120 1 0 $X=566680 $Y=597700
X86 3 11 61 19 INV1S $T=484840 613200 0 0 $X=484840 $Y=612820
X87 7 11 10 19 INV1S $T=491660 633360 1 0 $X=491660 $Y=627940
X88 9 11 1 19 INV1S $T=498480 603120 0 0 $X=498480 $Y=602740
X89 20 11 12 19 INV1S $T=516460 593040 0 0 $X=516460 $Y=592660
X90 24 11 17 19 INV1S $T=522660 593040 0 0 $X=522660 $Y=592660
X91 28 11 22 19 INV1S $T=529480 593040 0 0 $X=529480 $Y=592660
.ENDS
***************************************
.SUBCKT ND2 I1 O I2 GND VCC
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI22S A1 B1 O B2 GND A2 VCC
** N=10 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ND3 I3 GND I2 O VCC I1
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OR2 I2 I1 VCC GND O
** N=7 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT XOR2HS I1 I2 O VCC GND
** N=9 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MOAI1S B1 B2 GND A1 A2 O VCC
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OR3B2 I1 B1 VCC O B2 GND
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AO112 O C2 C1 VCC B1 GND A1
** N=10 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AO222 C1 C2 B2 B1 A1 A2 GND VCC O
** N=13 EP=9 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI12HS B2 B1 GND A1 VCC O
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AN2 I1 I2 GND VCC O
** N=7 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_21 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41
+ 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61
+ 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81
+ 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 98
** N=241 EP=96 IP=1011 FDC=0
X0 163 67 59 16 5 69 QDFFRBT $T=541880 492240 0 0 $X=541880 $Y=491860
X1 200 67 59 16 5 90 QDFFRBT $T=569160 492240 0 0 $X=569160 $Y=491860
X2 224 67 59 16 5 73 QDFFRBT $T=584040 512400 0 180 $X=570400 $Y=506980
X3 190 67 59 16 5 85 QDFFRBT $T=571020 522480 1 0 $X=571020 $Y=517060
X4 162 67 59 16 5 82 QDFFRBT $T=572880 502320 0 0 $X=572880 $Y=501940
X5 237 67 59 16 5 83 QDFFRBT $T=605120 502320 1 180 $X=591480 $Y=501940
X6 240 67 59 16 5 87 QDFFRBT $T=609460 502320 0 180 $X=595820 $Y=496900
X7 230 67 59 16 5 95 QDFFRBT $T=595820 522480 1 0 $X=595820 $Y=517060
X8 28 5 19 20 8 16 104 FA1S $T=476160 562800 0 0 $X=476160 $Y=562420
X9 109 5 30 26 28 16 117 FA1S $T=489800 562800 0 0 $X=489800 $Y=562420
X10 37 5 42 6 41 16 123 FA1S $T=496000 582960 0 0 $X=496000 $Y=582580
X11 124 5 26 111 125 16 130 FA1S $T=499100 532560 0 0 $X=499100 $Y=532180
X12 125 5 20 127 39 16 131 FA1S $T=499720 532560 1 0 $X=499720 $Y=527140
X13 138 5 51 46 141 16 148 FA1S $T=514600 552720 1 0 $X=514600 $Y=547300
X14 141 5 40 47 109 16 149 FA1S $T=515840 562800 0 0 $X=515840 $Y=562420
X15 142 5 47 134 124 16 135 FA1S $T=516460 532560 0 0 $X=516460 $Y=532180
X16 155 5 55 49 159 16 168 FA1S $T=526380 542640 1 0 $X=526380 $Y=537220
X17 156 5 46 150 142 16 133 FA1S $T=527000 512400 0 0 $X=527000 $Y=512020
X18 159 5 53 65 138 16 152 FA1S $T=539400 552720 0 180 $X=527620 $Y=547300
X19 166 5 157 158 170 16 206 FA1S $T=531340 572880 0 0 $X=531340 $Y=572500
X20 173 5 49 169 175 16 185 FA1S $T=540640 522480 1 0 $X=540640 $Y=517060
X21 175 5 65 171 156 16 193 FA1S $T=542500 512400 0 0 $X=542500 $Y=512020
X22 181 5 167 177 176 16 194 FA1S $T=546220 562800 0 0 $X=546220 $Y=562420
X23 191 5 180 182 181 16 202 FA1S $T=551180 562800 1 0 $X=551180 $Y=557380
X24 192 5 183 186 172 16 72 FA1S $T=551800 582960 1 0 $X=551800 $Y=577540
X25 208 5 166 194 209 16 217 FA1S $T=565440 562800 0 0 $X=565440 $Y=562420
X26 209 5 204 192 206 16 218 FA1S $T=565440 572880 1 0 $X=565440 $Y=567460
X27 211 5 205 191 210 16 225 FA1S $T=567300 552720 1 0 $X=567300 $Y=547300
X28 210 5 202 208 221 16 215 FA1S $T=570400 562800 1 0 $X=570400 $Y=557380
X29 219 5 214 213 79 16 226 FA1S $T=575980 582960 1 0 $X=575980 $Y=577540
X30 75 5 207 74 77 16 80 FA1S $T=575980 582960 0 0 $X=575980 $Y=582580
X31 221 5 217 220 236 16 229 FA1S $T=578460 562800 0 0 $X=578460 $Y=562420
X32 220 5 219 218 76 16 228 FA1S $T=578460 572880 1 0 $X=578460 $Y=567460
X33 233 5 226 81 84 16 91 FA1S $T=591480 582960 1 0 $X=591480 $Y=577540
X34 236 5 233 228 93 16 241 FA1S $T=603260 572880 1 0 $X=603260 $Y=567460
X35 12 5 13 101 16 NR2 $T=482360 562800 1 0 $X=482360 $Y=557380
X36 14 5 110 43 16 NR2 $T=503440 572880 0 0 $X=503440 $Y=572500
X37 45 5 112 48 16 NR2 $T=509640 572880 0 0 $X=509640 $Y=572500
X38 50 5 157 58 16 NR2 $T=523280 572880 1 0 $X=523280 $Y=567460
X39 50 5 167 57 16 NR2 $T=531340 562800 0 0 $X=531340 $Y=562420
X40 62 5 158 61 16 NR2 $T=536300 582960 1 180 $X=534440 $Y=582580
X41 56 5 170 63 16 NR2 $T=541260 582960 1 0 $X=541260 $Y=577540
X42 61 5 172 63 16 NR2 $T=542500 582960 0 0 $X=542500 $Y=582580
X43 66 5 176 63 16 NR2 $T=543120 572880 1 0 $X=543120 $Y=567460
X44 50 5 180 63 16 NR2 $T=546220 562800 1 0 $X=546220 $Y=557380
X45 62 5 177 56 16 NR2 $T=548080 582960 1 0 $X=548080 $Y=577540
X46 50 5 183 68 16 NR2 $T=548700 582960 0 0 $X=548700 $Y=582580
X47 62 5 182 66 16 NR2 $T=551800 572880 1 0 $X=551800 $Y=567460
X48 62 5 186 70 16 NR2 $T=554900 582960 0 0 $X=554900 $Y=582580
X49 62 5 205 50 16 NR2 $T=559240 552720 1 0 $X=559240 $Y=547300
X50 66 5 204 57 16 NR2 $T=559860 572880 1 0 $X=559860 $Y=567460
X51 61 5 207 57 16 NR2 $T=561100 582960 0 0 $X=561100 $Y=582580
X52 66 5 214 58 16 NR2 $T=567920 582960 1 0 $X=567920 $Y=577540
X53 56 5 213 57 16 NR2 $T=569780 582960 1 180 $X=567920 $Y=582580
X54 203 5 216 165 16 NR2 $T=568540 532560 1 0 $X=568540 $Y=527140
X55 15 9 102 16 5 103 HA1 $T=478640 512400 0 0 $X=478640 $Y=512020
X56 110 112 29 16 5 22 HA1 $T=499100 572880 1 180 $X=491040 $Y=572500
X57 113 108 115 16 5 128 HA1 $T=493520 512400 1 0 $X=493520 $Y=506980
X58 106 102 108 16 5 129 HA1 $T=502820 512400 0 0 $X=502820 $Y=512020
X59 136 115 144 16 5 146 HA1 $T=515840 512400 0 0 $X=515840 $Y=512020
X60 143 144 151 16 5 153 HA1 $T=522040 502320 0 0 $X=522040 $Y=501940
X61 184 151 187 16 5 196 HA1 $T=548700 512400 1 0 $X=548700 $Y=506980
X62 189 187 203 16 5 195 HA1 $T=556140 522480 1 0 $X=556140 $Y=517060
X63 17 5 101 16 INV1S $T=483600 532560 0 0 $X=483600 $Y=532180
X64 18 5 14 16 INV1S $T=483600 572880 0 0 $X=483600 $Y=572500
X65 27 5 9 16 INV1S $T=492900 502320 1 180 $X=491660 $Y=501940
X66 30 5 111 16 INV1S $T=494140 542640 1 0 $X=494140 $Y=537220
X67 32 5 99 16 INV1S $T=496620 552720 1 0 $X=496620 $Y=547300
X68 19 5 127 16 INV1S $T=508400 542640 0 180 $X=507160 $Y=537220
X69 131 5 106 16 INV1S $T=509020 522480 0 180 $X=507780 $Y=517060
X70 130 5 113 16 INV1S $T=510880 502320 1 180 $X=509640 $Y=501940
X71 49 5 50 16 INV1S $T=514600 582960 1 0 $X=514600 $Y=577540
X72 133 5 143 16 INV1S $T=516460 502320 0 0 $X=516460 $Y=501940
X73 135 5 136 16 INV1S $T=517080 522480 0 0 $X=517080 $Y=522100
X74 4 5 48 16 INV1S $T=517080 572880 0 0 $X=517080 $Y=572500
X75 46 5 56 16 INV1S $T=517700 582960 0 0 $X=517700 $Y=582580
X76 44 5 33 16 INV1S $T=518940 562800 1 0 $X=518940 $Y=557380
X77 40 5 134 16 INV1S $T=522040 542640 0 180 $X=520800 $Y=537220
X78 51 5 57 16 INV1S $T=525140 572880 0 0 $X=525140 $Y=572500
X79 51 5 150 16 INV1S $T=526380 522480 1 0 $X=526380 $Y=517060
X80 40 5 58 16 INV1S $T=526380 582960 0 0 $X=526380 $Y=582580
X81 55 5 169 16 INV1S $T=535680 522480 0 0 $X=535680 $Y=522100
X82 53 5 63 16 INV1S $T=536920 562800 0 0 $X=536920 $Y=562420
X83 55 5 62 16 INV1S $T=541880 562800 1 0 $X=541880 $Y=557380
X84 53 5 171 16 INV1S $T=542500 512400 1 0 $X=542500 $Y=506980
X85 65 5 66 16 INV1S $T=544980 582960 1 0 $X=544980 $Y=577540
X86 173 5 165 16 INV1S $T=547460 532560 1 0 $X=547460 $Y=527140
X87 185 5 189 16 INV1S $T=553660 522480 1 0 $X=553660 $Y=517060
X88 193 5 184 16 INV1S $T=561100 512400 1 0 $X=561100 $Y=506980
X89 165 5 178 16 INV1S $T=570400 532560 0 0 $X=570400 $Y=532180
X90 223 5 114 16 INV1S $T=586520 532560 1 0 $X=586520 $Y=527140
X91 155 188 12 16 5 ND2 $T=544360 532560 0 0 $X=544360 $Y=532180
X92 232 88 179 16 5 ND2 $T=595820 552720 0 0 $X=595820 $Y=552340
X93 231 230 179 16 5 ND2 $T=596440 532560 1 0 $X=596440 $Y=527140
X94 227 86 179 16 5 ND2 $T=596440 562800 1 0 $X=596440 $Y=557380
X95 235 237 179 16 5 ND2 $T=608840 532560 1 0 $X=608840 $Y=527140
X96 238 94 179 16 5 ND2 $T=608840 562800 1 0 $X=608840 $Y=557380
X97 239 240 179 16 5 ND2 $T=609460 532560 0 0 $X=609460 $Y=532180
X98 234 96 179 16 5 ND2 $T=614420 552720 1 0 $X=614420 $Y=547300
X99 3 99 2 9 16 10 5 AOI22S $T=480500 502320 0 0 $X=480500 $Y=501940
X100 3 99 11 15 16 100 5 AOI22S $T=481740 522480 1 0 $X=481740 $Y=517060
X101 27 107 1 27 16 114 5 AOI22S $T=491040 502320 1 0 $X=491040 $Y=496900
X102 3 99 118 106 16 105 5 AOI22S $T=494760 522480 1 180 $X=491040 $Y=522100
X103 103 107 21 31 16 114 5 AOI22S $T=493520 522480 1 0 $X=493520 $Y=517060
X104 3 99 116 113 16 121 5 AOI22S $T=499720 502320 0 0 $X=499720 $Y=501940
X105 128 107 119 130 16 114 5 AOI22S $T=507780 502320 1 0 $X=507780 $Y=496900
X106 129 107 120 131 16 114 5 AOI22S $T=507780 522480 0 0 $X=507780 $Y=522100
X107 3 99 139 136 16 132 5 AOI22S $T=520800 522480 0 180 $X=517080 $Y=517060
X108 146 107 147 135 16 114 5 AOI22S $T=525140 522480 0 0 $X=525140 $Y=522100
X109 3 99 160 143 16 140 5 AOI22S $T=530100 502320 0 180 $X=526380 $Y=496900
X110 153 107 161 133 16 114 5 AOI22S $T=534440 502320 0 0 $X=534440 $Y=501940
X111 165 178 179 99 16 101 5 AOI22S $T=550560 542640 0 180 $X=546840 $Y=537220
X112 3 99 199 184 16 174 5 AOI22S $T=555520 502320 0 180 $X=551800 $Y=496900
X113 196 107 198 193 16 114 5 AOI22S $T=558620 512400 0 0 $X=558620 $Y=512020
X114 216 215 227 35 16 114 5 AOI22S $T=575360 552720 1 180 $X=571640 $Y=552340
X115 212 78 222 35 16 114 5 AOI22S $T=582800 542640 1 0 $X=582800 $Y=537220
X116 216 211 234 35 16 114 5 AOI22S $T=588380 552720 0 180 $X=584660 $Y=547300
X117 216 225 232 35 16 114 5 AOI22S $T=595200 542640 0 0 $X=595200 $Y=542260
X118 216 89 231 35 16 114 5 AOI22S $T=595820 532560 0 0 $X=595820 $Y=532180
X119 216 92 235 35 16 114 5 AOI22S $T=608220 542640 0 180 $X=604500 $Y=537220
X120 216 229 238 35 16 114 5 AOI22S $T=607600 552720 0 0 $X=607600 $Y=552340
X121 216 241 239 35 16 114 5 AOI22S $T=608220 542640 0 0 $X=608220 $Y=542260
X122 222 16 188 224 5 179 ND3 $T=582800 532560 0 0 $X=582800 $Y=532180
X123 178 64 5 16 223 OR2 $T=577220 532560 1 0 $X=577220 $Y=527140
X124 18 23 10 5 16 XOR2HS $T=478640 552720 1 0 $X=478640 $Y=547300
X125 4 7 100 5 16 XOR2HS $T=480500 532560 1 0 $X=480500 $Y=527140
X126 20 19 105 5 16 XOR2HS $T=484840 542640 1 0 $X=484840 $Y=537220
X127 26 30 121 5 16 XOR2HS $T=498480 542640 1 0 $X=498480 $Y=537220
X128 47 40 132 5 16 XOR2HS $T=511500 542640 1 0 $X=511500 $Y=537220
X129 46 51 140 5 16 XOR2HS $T=516460 502320 1 0 $X=516460 $Y=496900
X130 49 55 154 5 16 XOR2HS $T=526380 532560 1 0 $X=526380 $Y=527140
X131 65 53 174 5 16 XOR2HS $T=541880 502320 1 0 $X=541880 $Y=496900
X132 203 178 212 5 16 XOR2HS $T=569160 542640 1 0 $X=569160 $Y=537220
X133 71 35 16 185 32 201 5 MOAI1S $T=564820 542640 1 180 $X=561100 $Y=542260
X134 126 119 5 36 116 16 OR3B2 $T=503440 502320 0 180 $X=499720 $Y=496900
X135 122 120 5 38 118 16 OR3B2 $T=503440 522480 1 180 $X=499720 $Y=522100
X136 164 147 5 162 139 16 OR3B2 $T=536920 522480 0 180 $X=533200 $Y=517060
X137 137 161 5 163 160 16 OR3B2 $T=538160 502320 0 180 $X=534440 $Y=496900
X138 145 198 5 200 199 16 OR3B2 $T=562960 502320 0 180 $X=559240 $Y=496900
X139 190 12 168 5 197 16 201 AO112 $T=555520 532560 0 0 $X=555520 $Y=532180
X140 104 12 33 30 34 35 16 5 122 AO222 $T=496000 552720 0 0 $X=496000 $Y=552340
X141 117 12 33 40 123 35 16 5 126 AO222 $T=499720 562800 1 0 $X=499720 $Y=557380
X142 148 12 33 53 52 35 16 5 137 AO222 $T=524520 542640 1 180 $X=518320 $Y=542260
X143 152 12 33 55 54 35 16 5 145 AO222 $T=528860 552720 1 180 $X=522660 $Y=552340
X144 149 12 33 51 60 35 16 5 164 AO222 $T=529480 562800 1 0 $X=529480 $Y=557380
X145 3 154 114 195 107 185 16 5 197 AO222 $T=555520 532560 1 0 $X=555520 $Y=527140
X146 64 165 16 17 5 107 OAI12HS $T=537540 532560 1 180 $X=533820 $Y=532180
X147 18 23 16 5 25 AN2 $T=486080 572880 1 0 $X=486080 $Y=567460
.ENDS
***************************************
.SUBCKT TIE1 O VCC GND
** N=5 EP=3 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_22 3 4 5 10
** N=10 EP=4 IP=4 FDC=0
X0 3 5 4 TIE1 $T=672080 391440 0 0 $X=672080 $Y=391060
.ENDS
***************************************
.SUBCKT BUF2 I O GND VCC
** N=6 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_23 3 5 12 13 26
** N=26 EP=5 IP=5 FDC=0
X0 3 5 12 13 BUF2 $T=557380 341040 1 0 $X=557380 $Y=335620
.ENDS
***************************************
.SUBCKT ICV_24 5 6 7 8 9 10 25
** N=35 EP=7 IP=16 FDC=0
X0 5 6 7 7 7 8 7 YA2GSC $T=611160 0 0 0 $X=613070 $Y=0
X1 9 6 7 7 7 10 7 YA2GSC $T=669680 0 0 0 $X=671590 $Y=0
.ENDS
***************************************
.SUBCKT ICV_25 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=18 FDC=0
X0 1 3 1 1 2 XMC $T=384160 1110080 0 180 $X=351970 $Y=875100
X1 1 5 1 1 4 XMC $T=433680 1110080 0 180 $X=401490 $Y=875100
X2 1 7 1 1 6 XMC $T=483200 1110080 0 180 $X=451010 $Y=875100
.ENDS
***************************************
.SUBCKT BUF12CK I GND VCC O
** N=6 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_26 1 2 7 8 9 11
** N=11 EP=6 IP=10 FDC=0
X0 9 7 8 2 BUF12CK $T=345960 764400 0 0 $X=345960 $Y=764020
X1 9 7 8 1 BUF12CK $T=345960 774480 1 0 $X=345960 $Y=769060
.ENDS
***************************************
.SUBCKT ICV_27 1 2 3 4 5 6 7 8 13
** N=13 EP=9 IP=14 FDC=0
X0 1 2 3 8 7 5 QDFFRBN $T=372620 663600 0 0 $X=372620 $Y=663220
X1 4 2 3 8 7 6 QDFFRBN $T=388120 673680 0 0 $X=388120 $Y=673300
.ENDS
***************************************
.SUBCKT ICV_28 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 22
** N=22 EP=17 IP=39 FDC=0
X0 2 3 4 16 1 6 QDFFRBN $T=373240 653520 0 0 $X=373240 $Y=653140
X1 5 3 4 16 1 10 QDFFRBN $T=386260 633360 0 0 $X=386260 $Y=632980
X2 7 3 4 16 1 11 QDFFRBN $T=390600 603120 1 0 $X=390600 $Y=597700
X3 8 3 4 16 1 9 QDFFRBN $T=394940 653520 1 0 $X=394940 $Y=648100
X4 13 16 14 15 1 NR2 $T=468100 593040 0 0 $X=468100 $Y=592660
X5 11 16 12 1 INV1S $T=463140 603120 1 0 $X=463140 $Y=597700
.ENDS
***************************************
.SUBCKT OAI112HS C2 C1 GND B1 O A1 VCC
** N=9 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OA222 A2 A1 B2 B1 C2 C1 GND VCC O
** N=13 EP=9 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT XNR2HS I1 I2 O VCC GND
** N=9 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI12HS B2 B1 VCC A1 GND O
** N=8 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NR3 I1 VCC I2 I3 O GND
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MAOI1 B1 B2 A1 A2 VCC GND O
** N=10 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_29 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 48 49 50 51 53 55 56 57 58 61
** N=91 EP=56 IP=343 FDC=0
X0 62 3 5 44 46 2 QDFFRBT $T=380060 492240 1 180 $X=366420 $Y=491860
X1 68 3 5 44 46 11 QDFFRBT $T=427180 502320 1 180 $X=413540 $Y=501940
X2 19 3 5 44 46 14 QDFFRBT $T=451980 492240 1 180 $X=438340 $Y=491860
X3 25 3 5 44 46 17 QDFFRBT $T=457560 502320 0 180 $X=443920 $Y=496900
X4 1 3 5 46 44 6 QDFFRBN $T=361460 502320 1 0 $X=361460 $Y=496900
X5 4 3 5 46 44 12 QDFFRBN $T=368900 512400 1 0 $X=368900 $Y=506980
X6 7 3 5 46 44 13 QDFFRBN $T=394320 492240 0 0 $X=394320 $Y=491860
X7 8 3 5 46 44 26 QDFFRBN $T=397420 512400 0 0 $X=397420 $Y=512020
X8 9 3 5 46 44 10 QDFFRBN $T=398040 502320 1 0 $X=398040 $Y=496900
X9 63 3 5 46 44 66 QDFFRBN $T=417880 542640 0 0 $X=417880 $Y=542260
X10 64 3 5 46 44 65 QDFFRBN $T=422840 562800 0 0 $X=422840 $Y=562420
X11 71 3 5 46 44 76 QDFFRBN $T=442680 532560 1 0 $X=442680 $Y=527140
X12 21 46 24 12 22 44 75 FA1S $T=464380 562800 1 180 $X=452600 $Y=562420
X13 39 46 12 78 90 44 40 FA1S $T=468100 522480 0 0 $X=468100 $Y=522100
X14 55 46 57 58 56 44 43 FA1S $T=486080 582960 0 180 $X=474300 $Y=577540
X15 30 46 86 16 44 NR2 $T=468100 572880 1 180 $X=466240 $Y=572500
X16 45 46 85 49 44 NR2 $T=474920 572880 0 0 $X=474920 $Y=572500
X17 66 46 67 44 INV1S $T=440820 542640 0 0 $X=440820 $Y=542260
X18 15 46 72 44 INV1S $T=442680 572880 0 0 $X=442680 $Y=572500
X19 65 46 70 44 INV1S $T=443300 532560 0 0 $X=443300 $Y=532180
X20 76 46 73 44 INV1S $T=450120 542640 1 180 $X=448880 $Y=542260
X21 24 46 78 44 INV1S $T=460660 522480 1 180 $X=459420 $Y=522100
X22 6 46 88 44 INV1S $T=465620 522480 1 0 $X=465620 $Y=517060
X23 41 46 83 44 INV1S $T=469960 512400 0 180 $X=468720 $Y=506980
X24 40 46 51 44 INV1S $T=473060 512400 0 0 $X=473060 $Y=512020
X25 87 46 53 44 INV1S $T=475540 532560 0 0 $X=475540 $Y=532180
X26 80 46 33 44 INV1S $T=479260 542640 1 0 $X=479260 $Y=537220
X27 16 77 72 44 46 ND2 $T=451360 572880 0 180 $X=449500 $Y=567460
X28 41 90 88 44 46 ND2 $T=473680 522480 1 0 $X=473680 $Y=517060
X29 18 44 16 74 46 15 ND3 $T=444540 562800 1 180 $X=442060 $Y=562420
X30 65 44 67 20 46 76 ND3 $T=455080 532560 0 0 $X=455080 $Y=532180
X31 76 44 70 23 46 67 ND3 $T=456940 542640 0 0 $X=456940 $Y=542260
X32 65 44 73 80 46 67 ND3 $T=460040 552720 0 180 $X=457560 $Y=547300
X33 76 44 70 87 46 66 ND3 $T=466240 532560 0 0 $X=466240 $Y=532180
X34 65 44 73 31 46 66 ND3 $T=466860 552720 1 0 $X=466860 $Y=547300
X35 66 44 73 50 46 70 ND3 $T=472440 542640 1 0 $X=472440 $Y=537220
X36 69 16 44 69 67 63 46 MOAI1S $T=443920 552720 0 180 $X=440200 $Y=547300
X37 69 15 44 69 70 64 46 MOAI1S $T=445780 552720 1 180 $X=442060 $Y=552340
X38 69 18 44 69 73 71 46 MOAI1S $T=452600 552720 0 180 $X=448880 $Y=547300
X39 84 74 44 77 20 69 46 MOAI1S $T=458180 552720 1 180 $X=454460 $Y=552340
X40 81 27 46 62 37 44 OR3B2 $T=464380 502320 1 0 $X=464380 $Y=496900
X41 82 29 46 68 38 44 OR3B2 $T=465000 512400 0 0 $X=465000 $Y=512020
X42 75 28 32 34 36 33 44 46 82 AO222 $T=466860 562800 1 0 $X=466860 $Y=557380
X43 42 28 32 24 85 33 44 46 81 AO222 $T=474300 542640 1 180 $X=468100 $Y=542260
X44 23 77 44 91 84 48 46 OAI112HS $T=472440 552720 0 0 $X=472440 $Y=552340
X45 80 86 87 79 31 89 44 46 91 OA222 $T=469340 562800 0 0 $X=469340 $Y=562420
X46 83 6 35 46 44 XNR2HS $T=466860 502320 0 0 $X=466860 $Y=501940
X47 18 15 46 30 44 89 AOI12HS $T=465000 582960 1 0 $X=465000 $Y=577540
X48 65 46 76 66 28 44 NR3 $T=468100 542640 0 180 $X=465000 $Y=537220
X49 16 18 16 72 46 44 79 MAOI1 $T=453220 572880 0 0 $X=453220 $Y=572500
.ENDS
***************************************
.SUBCKT ICV_30
** N=8 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_31
** N=9 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_32 1 2 3 4 5 6 7
** N=7 EP=7 IP=16 FDC=0
X0 1 2 3 3 3 4 3 YA2GSC $T=377080 0 0 0 $X=378990 $Y=0
X1 5 2 3 3 3 6 3 YA2GSC $T=435600 0 0 0 $X=437510 $Y=0
.ENDS
***************************************
.SUBCKT ICV_33 1 2 3 4 5 6 7
** N=7 EP=7 IP=12 FDC=0
X0 1 3 1 1 2 XMC $T=1110080 -334640 0 90 $X=875100 $Y=-332790
X1 4 6 4 4 5 XMC $T=1110080 -285120 0 90 $X=875100 $Y=-283270
.ENDS
***************************************
.SUBCKT ICV_34
** N=10 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT BUF3 I VCC GND O
** N=6 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_35 1 5 6 7 9
** N=9 EP=5 IP=5 FDC=0
X0 7 6 5 1 BUF3 $T=347200 673680 0 0 $X=347200 $Y=673300
.ENDS
***************************************
.SUBCKT ICV_36
** N=8 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_37
** N=8 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_38
** N=8 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_39
** N=11 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_40 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=16 FDC=0
X0 1 2 3 3 3 4 3 YA2GSC $T=0 -318560 0 270 $X=0 $Y=-351430
X1 5 2 6 6 6 7 3 YA2GSC $T=0 -260030 0 270 $X=0 $Y=-292900
.ENDS
***************************************
.SUBCKT ICV_41
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_42 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=18 FDC=0
X0 2 5 2 2 1 XMC $T=0 764370 0 270 $X=0 $Y=732180
X1 2 6 2 2 3 XMC $T=0 812440 0 270 $X=0 $Y=780250
X2 2 7 2 2 4 XMC $T=0 860510 0 270 $X=0 $Y=828320
.ENDS
***************************************
.SUBCKT ICV_43 1 2 3 4
** N=4 EP=4 IP=6 FDC=0
X0 2 3 2 2 1 XMC $T=0 716300 0 270 $X=0 $Y=684110
.ENDS
***************************************
.SUBCKT ICV_44 1 2 3 4 5 6
** N=6 EP=6 IP=12 FDC=0
X0 1 3 1 1 2 XMC $T=0 620160 0 270 $X=0 $Y=587970
X1 1 5 1 1 4 XMC $T=0 668230 0 270 $X=0 $Y=636040
.ENDS
***************************************
.SUBCKT ICV_45 1 2 3 4
** N=14 EP=4 IP=6 FDC=0
X0 2 3 2 2 1 XMC $T=0 475950 0 270 $X=0 $Y=443760
.ENDS
***************************************
.SUBCKT ICV_46 1 2 3 4
** N=4 EP=4 IP=6 FDC=0
X0 2 3 2 2 1 XMC $T=0 427880 0 270 $X=0 $Y=395690
.ENDS
***************************************
.SUBCKT ICV_47 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=18 FDC=0
X0 2 5 2 2 1 XMC $T=0 283670 0 270 $X=0 $Y=251480
X1 2 6 2 2 3 XMC $T=0 331740 0 270 $X=0 $Y=299550
X2 2 7 2 2 4 XMC $T=0 379810 0 270 $X=0 $Y=347620
.ENDS
***************************************
.SUBCKT ICV_48
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT CHIP data_o[14] data_o[15] data_o[13] data_o[12] data_o[11] data_o[10] data_o[8] data_o[9] data_a_i[4] data_a_i[3] GND VCC data_o[7] data_o[6] data_a_i[0] data_a_i[1] data_a_i[2] data_o[4] data_o[5] inst_i[0]
+ inst_i[1] inst_i[2] data_o[2] data_o[3] reset_n_i clk_p_i data_o[1] data_o[0] data_b_i[5] data_b_i[6] data_b_i[7] data_b_i[4] data_b_i[2] data_b_i[3] data_b_i[1] data_b_i[0] data_a_i[5] data_a_i[6] data_a_i[7]
** N=213 EP=39 IP=652 FDC=0
X1 1 2 3 4 data_o[14] data_o[15] 213 ICV_2 $T=0 0 0 0 $X=845870 $Y=732200
X2 1 2 7 data_o[13] 213 ICV_3 $T=0 0 0 0 $X=845870 $Y=662600
X3 data_o[12] 1 2 161 213 ICV_4 $T=0 0 0 0 $X=845870 $Y=588000
X4 1 2 11 data_o[11] 213 ICV_5 $T=0 0 0 0 $X=845870 $Y=448100
X5 1 13 14 data_o[10] 213 ICV_6 $T=0 0 0 0 $X=845870 $Y=378000
X6 1 13 16 17 data_o[8] data_o[9] 213 ICV_7 $T=0 0 0 0 $X=845870 $Y=235000
X8 2 24 data_a_i[4] 98 data_a_i[3] 213 ICV_9 $T=0 0 0 90 $X=729000 $Y=875100
X13 2 13 VCC GND 213 ICV_14 $T=0 0 0 0 $X=729000 $Y=378000
X15 data_o[7] 1 25 13 100 data_o[6] 99 213 ICV_16 $T=0 0 0 90 $X=729000 $Y=0
X16 2 105 data_a_i[0] 106 data_a_i[1] 107 data_a_i[2] 213 ICV_17 $T=0 0 0 0 $X=481400 $Y=875100
X18 39 108 68 168 106 107 42 2 105 109 98 110 4 199 3 24 111 VCC GND 213 ICV_19 $T=0 0 0 0 $X=481400 $Y=662600
X19 36 37 39 52 112 55 113 201 42 129 VCC 125 116 114 115 35 117 200 GND 118
+ 120 124 119 108 121 122 123 109 131 128 126 203 127 202 130 132 133 138 134 135
+ 137 139 136 140 141 161 168 68 142 7 143 144 145 213
+ ICV_20 $T=0 0 0 0 $X=478640 $Y=587620
X20 47 45 43 46 VCC 53 108 186 40 49 176 51 50 52 174 GND 48 41 39 38
+ 175 184 42 187 113 172 44 54 109 177 181 183 188 182 170 115 173 179 199 114
+ 116 117 185 36 156 118 120 167 122 171 200 169 201 178 119 128 123 68 121 125
+ 126 127 180 157 131 168 124 146 129 202 132 16 133 134 135 130 136 203 137 138
+ 147 14 140 100 141 11 110 139 99 142 145 143 144 17 111 213
+ ICV_21 $T=0 0 0 0 $X=476160 $Y=448100
X21 1 GND VCC 213 ICV_22 $T=0 0 0 0 $X=481400 $Y=378000
X22 2 25 GND VCC 213 ICV_23 $T=0 0 0 0 $X=481400 $Y=235000
X23 data_o[4] 1 25 147 data_o[5] 146 213 ICV_24 $T=0 0 0 0 $X=481400 $Y=0
X24 2 152 inst_i[0] 153 inst_i[1] 154 inst_i[2] 213 ICV_25 $T=0 0 0 0 $X=351970 $Y=875100
X25 168 155 GND VCC 65 213 ICV_26 $T=0 0 0 0 $X=345960 $Y=732200
X26 67 155 68 66 156 167 GND VCC 213 ICV_27 $T=0 0 0 0 $X=352000 $Y=662600
X27 GND 70 155 68 69 157 193 81 118 113 38 37 153 158 154 VCC 213 ICV_28 $T=0 0 0 0 $X=352000 $Y=588000
X28 72 75 155 71 68 41 83 73 82 171 74 46 169 159 153 152 160 154 173 180
+ 186 187 181 108 170 178 47 51 175 158 185 183 182 39 172 184 45 176 179 177
+ 42 49 188 GND 36 VCC 50 52 48 174 43 53 112 55 54 213
+ ICV_29 $T=0 0 0 0 $X=352000 $Y=448100
X31 data_o[2] 1 25 159 data_o[3] 160 213 ICV_32 $T=0 0 0 0 $X=352000 $Y=0
X32 2 68 reset_n_i 80 65 clk_p_i 213 ICV_33 $T=0 0 0 90 $X=235000 $Y=875100
X34 80 GND VCC 2 213 ICV_35 $T=0 0 0 0 $X=235000 $Y=662600
X39 data_o[1] 1 25 74 data_o[0] 80 75 213 ICV_40 $T=0 0 0 90 $X=235000 $Y=0
X41 67 80 70 66 data_b_i[5] data_b_i[6] data_b_i[7] 213 ICV_42 $T=0 0 0 0 $X=0 $Y=732180
X42 81 80 data_b_i[4] 213 ICV_43 $T=0 0 0 0 $X=0 $Y=662600
X43 80 193 data_b_i[2] 69 data_b_i[3] 213 ICV_44 $T=0 0 0 0 $X=0 $Y=587970
X44 71 80 data_b_i[1] 213 ICV_45 $T=0 0 0 0 $X=0 $Y=443760
X45 72 80 data_b_i[0] 213 ICV_46 $T=0 0 0 0 $X=0 $Y=378000
X46 82 80 83 73 data_a_i[5] data_a_i[6] data_a_i[7] 213 ICV_47 $T=0 0 0 0 $X=0 $Y=235000
.ENDS
***************************************
